module rain

enum Token {

}

