module rain

enum Tokens {
	
}

